module seg (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n // Asynchronous reset active low
	
);

endmodule