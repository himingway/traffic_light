module traffic_light (
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	output[1:0] light_control
);

endmodule